----------------------------------------------------------------------------------
-- Company: 
-- Engineer: 
-- 
-- Create Date:    14:31:22 12/07/2012 
-- Design Name: 
-- Module Name:    muxI - Behavioral 
-- Project Name: 
-- Target Devices: 
-- Tool versions: 
-- Description: 
--
-- Dependencies: 
--
-- Revision: 
-- Revision 0.01 - File Created
-- Additional Comments: 
--
----------------------------------------------------------------------------------
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

-- Uncomment the following library declaration if using
-- arithmetic functions with Signed or Unsigned values
--use IEEE.NUMERIC_STD.ALL;

-- Uncomment the following library declaration if instantiating
-- any Xilinx primitives in this code.
--library UNISIM;
--use UNISIM.VComponents.all;

entity muxI is
    Port ( inst1 : in  STD_LOGIC_VECTOR (15 downto 0);
           inst2 : in  STD_LOGIC_VECTOR (15 downto 0);
           s : in  STD_LOGIC;
           instout : out  STD_LOGIC_VECTOR (15 downto 0));
end muxI;

architecture Behavioral of muxI is

begin
process(s) begin
	if (s='0') then
		instout<=inst1;
	else
		instout<=inst2;
	end if;	
end process;		


end Behavioral;

